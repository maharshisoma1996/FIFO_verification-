
`define data_width 8
`define d_out_width 8
`define fifo_depth 32


