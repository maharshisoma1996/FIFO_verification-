
`include "default_widths.sv"

`include "interface.sv"
`include "transcation.sv"
`include "generator.sv"
`include "driver.sv"

`include "monitor.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include"ram.txt"
`include"syn_fifo.txt"
